/*
Author: Sajeed Mohammad Shahriat
Affiliation: Rochester Institute of Technology
All rights reserved
This files can be reused and modified given that this copyright notice is not removed
*/

module comparator (
	a,
	b,
	a_less_b,
	a_equal_b,
	a_greater_b

); //end of port list

//---------------------------input ports-----------------------------


//---------------------------output ports----------------------------


//-----------------------input port data type------------------------


//-----------------------output port data type-----------------------


//---------------------------RTL design------------------------------

endmodule 
