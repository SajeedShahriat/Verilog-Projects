/*
Author: Sajeed Mohammad Shahriat
Affiliation: Rochester Institute of Technology
All rights reserved
This files can be reused and modified given that this copyright notice is not removed
*/

module (



); //end of port list

//---------------------------input ports-----------------------------


//---------------------------output ports----------------------------


//-----------------------input port data type------------------------


//-----------------------output port data type-----------------------


//---------------------------RTL design------------------------------

endmodule 
